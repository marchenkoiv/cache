`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 13.04.2023 00:30:08
// Design Name: 
// Module Name: tb_muu
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_if();

    reg areset = 'b0;
    reg sys_clk = 'b0;
    reg c_clk = 'b0;
    reg ram_clk = 'b0;
    reg [15:0] addr;
    reg wr = 'b0;
    reg rd = 'b0;
    reg [31:0] wdata;
    reg [3:0] bval;
    
    reg [7:0] rrdata;
    reg rack = 'b0;
    
    wire [31:0] rdata;
    wire ack;
    
    wire [12:0] raddr;
    wire rnw;
    wire [7:0]rwdata;
    wire avalid;
    
    
    
    cache dut(

    sys_clk,
    c_clk,
    ram_clk,
    addr,
    wr,
    rd,
    wdata,
    bval,
    areset,
    rrdata,
    rack,
    rdata,
    ack,
    raddr,
    rnw,
    rwdata,
    avalid
    );
    
    always #2 sys_clk <= ~sys_clk;
    always #7 c_clk <= ~c_clk;
    always #23 ram_clk <= ~ram_clk;
    
    initial #100 begin : test
        #10
        
        areset <= 'b1;
        #20
        areset <= 'b0;
        $display("test begin");
        
//                @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        rd = 'b0;
//        wr = 'b1;
//        addr = 'b0;
//        bval = 'b0001;
//        @(posedge sys_clk);
//        wr = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        rd = 'b0;
//        wr = 'b1;
//        addr = 'b01_000000_000;
//        bval = 'b0001;
//        @(posedge sys_clk);
//        wr = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160
         
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b10_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160       
   
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b11_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160     
        
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        rd = 'b0;
//        wr = 'b1;
//        addr = 'b100_000000_000;
//        bval = 'b0001;
//        @(posedge sys_clk);
//        wr = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160
 
//        @(posedge sys_clk);
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b101_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160 
 
//        @(posedge sys_clk);
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b110_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160 
        
//        @(posedge sys_clk);
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b111_000000_000;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160 
        
//        @(posedge sys_clk);
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b1000_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        @(posedge ram_clk);
//        rack = 'b0;
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rrdata = $urandom%63;
//        rack = 'b1;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #160
        
//        @(posedge sys_clk);
//        wr = 'b1;
//        rd = 'b0;
//        addr = 'b1001_000000_100;
//        bval = 'b0001;
//        @(posedge sys_clk);
//        wr = 'b0;
//        addr = 'b0;
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        @(posedge ram_clk);
//        rack = 'b0;
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge c_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b1;
//        rrdata = $urandom%63;
//        @(posedge ram_clk);
//        rack = 'b0;
//        rrdata = 'b0;
//        #200
        
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        wr = 'b0;
//        rd = 'b1;
//        addr = 'b10_000000_100;
//        bval = 'b0000;
//        @(posedge sys_clk);
//        rd = 'b0;
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
        
//        @(posedge sys_clk);
//        wdata = 'b10101010101;
//        //RData = 'b11111111111;
//        wr = 'b1;
//        rd = 'b0;
//        addr = 'b10_000000_100;
//        bval = 'b0001;
//        @(posedge sys_clk);
//        rd = 'b0;
//        wr = 'b0; 
//        addr = 'b0;
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        @(posedge ram_clk);
//        #50
        
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        rd = 'b0;
        wr = 'b1;
        addr = 'b0;
        bval = 'b0001;
        @(posedge sys_clk);
        wr = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        rd = 'b0;
        wr = 'b1;
        addr = 'b01_000000_000;
        bval = 'b0001;
        @(posedge sys_clk);
        wr = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160
         
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        wr = 'b0;
        rd = 'b1;
        addr = 'b10_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160       
   
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        wr = 'b0;
        rd = 'b1;
        addr = 'b11_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160     
        
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        rd = 'b0;
        wr = 'b1;
        addr = 'b100_000000_000;
        bval = 'b0001;
        @(posedge sys_clk);
        wr = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160
 
        @(posedge sys_clk);
        wr = 'b0;
        rd = 'b1;
        addr = 'b101_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160 
 
        @(posedge sys_clk);
        wr = 'b0;
        rd = 'b1;
        addr = 'b110_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160 
        
        @(posedge sys_clk);
        wr = 'b0;
        rd = 'b1;
        addr = 'b111_000000_000;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160 
        
        @(posedge sys_clk);
        wr = 'b0;
        rd = 'b1;
        addr = 'b1000_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        @(posedge ram_clk);
        rack = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rrdata = $urandom%63;
        rack = 'b1;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #160
        
        @(posedge sys_clk);
        wr = 'b1;
        rd = 'b0;
        addr = 'b1001_000000_100;
        bval = 'b0001;
        @(posedge sys_clk);
        wr = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        @(posedge ram_clk);
        rack = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b1;
        rrdata = $urandom%63;
        @(posedge ram_clk);
        rack = 'b0;
        rrdata = 'b0;
        #200
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        wr = 'b0;
        rd = 'b1;
        addr = 'b10_000000_100;
        bval = 'b0000;
        @(posedge sys_clk);
        rd = 'b0;
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
        
        @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        wr = 'b1;
        rd = 'b0;
        addr = 'b10_000000_100;
        bval = 'b0001;
        @(posedge sys_clk);
        rd = 'b0;
        wr = 'b0; 
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);
                @(posedge sys_clk);
        wdata = 'b10101010101;
        //RData = 'b11111111111;
        wr = 'b1;
        rd = 'b0;
        addr = 'b10_000000_100;
        bval = 'b0010;
        @(posedge sys_clk);
        rd = 'b0;
        wr = 'b0; 
        addr = 'b0;
        @(posedge ram_clk);
        @(posedge ram_clk);
        @(posedge ram_clk);

        #50
        

        
        $display("test end");
        $finish;
    end : test
endmodule
